module alu (
    input  [31:0] a,
    input  [31:0] b,
    input  [2:0]  alu_ctrl,
    output reg [31:0] result,
    output        zero
);

    wire signed [31:0] a_signed;
    wire signed [31:0] b_signed;

    assign a_signed = a;
    assign b_signed = b;

    always @(*) begin
        case (alu_ctrl)
            3'b000: result = a + b;                       // ADD
            3'b001: result = a - b;                       // SUB
            3'b010: result = a & b;                       // AND
            3'b011: result = a | b;                       // OR
            3'b100: result = a ^ b;                       // XOR
            3'b101: result = (a_signed < b_signed) ? 32'd1 : 32'd0; // SLT
            default: result = 32'd0;
        endcase
    end

    assign zero = (result == 32'd0);

endmodule

